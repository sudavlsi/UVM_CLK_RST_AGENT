class clk_rst_cfg extends uvm_object;
	`uvm_object_utils(clk_rst_cfg)

	function new();

	endfunction

endclass
