interface uvm_clk_rst_intf#( BIT_WIDTH = 1 , NUM_STAGES = 2 );
   logic clk, rstN;


endinterface
