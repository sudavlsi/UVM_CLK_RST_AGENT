package clk_rst_pkg;
	`include "clk_rst_cfg.sv"
	`include "clk_rst_agent.sv"
endpackage
